package env_pkg;

  import agent_pkg::*;

  `include "fifo_sco.sv"
  `include "fifo_env.sv"

endpackage