package agent_pkg;

    `include "fifo_trans.sv"
    `include "fifo_driver.sv"
    `include "fifo_monitor.sv"
    `include "fifo_generator.sv"
    

endpackage